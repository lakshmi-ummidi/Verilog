/********************************************************************************************

Filename    :	   half_adder.v   

Description :      Half adder Design using dataflow model

Author Name :      Lakshmi Ummidi

Version     :      1.0
*********************************************************************************************/
  
module half_adder(a, b, sum,carry);

	input a,b;
	output sum,carry;
   //Understand the Data-flow abstraction
   assign sum   = a ^ b;
   assign carry = a & b;

endmodule
	
	
	
	

	
	
